package tb_pkg;
// import uvm_pkg::*;
 // `include "uvm_macros.svh"
`include "packet.sv"
`include "transaction.sv"
`include "axi_sequence.sv"
`include "apb_sequence.sv"
`include "axi_driver.sv"
`include "apb_driver.sv"
`include "axi_monitor.sv"
`include "apb_monitor.sv"
`include "scoreboard.sv"
`include "axi_agent.sv"
`include "apb_agent.sv"
`include "environment.sv"
//`include "test_collection.sv"
//`include "test.sv"


endpackage
